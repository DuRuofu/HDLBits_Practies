module top_module( input in, output out );
	assign out =!in;
    //or 
    //assign out =~in;
endmodule
